`define BITWIDTH        8
`define FULLBITWIDTH    32
`define ADDR_WIDTH      18
`define MODE_ADDR_WIDTH 2


`define AXI_DONE_ADDR           40'h04_0004_0000
`define AXI_START_ADDR          40'h04_0008_0000
`define AXI_TRANSFER_MASK       16'h04_0

`define AXI_DATA_WIDTH              32